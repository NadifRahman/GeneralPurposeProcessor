library verilog;
use verilog.vl_types.all;
entity GPP_vlg_vec_tst is
end GPP_vlg_vec_tst;
