library verilog;
use verilog.vl_types.all;
entity mealy10circuit_vlg_vec_tst is
end mealy10circuit_vlg_vec_tst;
