library verilog;
use verilog.vl_types.all;
entity dec3to8_vlg_vec_tst is
end dec3to8_vlg_vec_tst;
