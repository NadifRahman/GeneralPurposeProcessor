library verilog;
use verilog.vl_types.all;
entity latch1_vlg_vec_tst is
end latch1_vlg_vec_tst;
