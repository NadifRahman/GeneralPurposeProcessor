library verilog;
use verilog.vl_types.all;
entity modifieddec4to16_vlg_vec_tst is
end modifieddec4to16_vlg_vec_tst;
